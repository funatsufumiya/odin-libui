module main

import libui

fn main() {
	println("hello")
}